`define WRITE 2'b00
`define JUMP 2'b01
`define BOTH 2'b10

module rob#(parameter ROB_WIDTH = 4)
           ();
    
endmodule //rob
