module decoder(
  input wire clk_in,
  input wire rdy_in,
  input [31:0] instruction
);


    
endmodule //decoder