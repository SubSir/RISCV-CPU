module if (input wire [7:0] mem_din,
           input wire from_lsb,
           output reg [7:0] mem_dout,
           output reg [31:0] mem_a,
           output reg mem_wr,
           );

endmodule //if
